module priority_deshiphrator (
    input [7:0] num,
    output reg [2:0] ub
);

    reg [2:0] a [7:0];
    reg [2:0] c [3:0];
    reg [2:0] d [1:0];

    always @(*) begin
        a[0] = (num[0]) ? 3'b000 : 3'b000;
        a[1] = (num[1]) ? 3'b001 : 3'b000;
        a[2] = (num[2]) ? 3'b010 : 3'b000;
        a[3] = (num[3]) ? 3'b011 : 3'b000;
        a[4] = (num[4]) ? 3'b100 : 3'b000;
        a[5] = (num[5]) ? 3'b101 : 3'b000;
        a[6] = (num[6]) ? 3'b110 : 3'b000;
        a[7] = (num[7]) ? 3'b111 : 3'b000;

        c[0] = (a[1] >= a[0]) ? a[1] : a[0];
        c[1] = (a[3] >= a[2]) ? a[3] : a[2];
        c[2] = (a[5] >= a[4]) ? a[5] : a[4];
        c[3] = (a[7] >= a[6]) ? a[7] : a[6];

        d[0] = (c[1] >= c[0]) ? c[1] : c[0];
        d[1] = (c[3] >= c[2]) ? c[3] : c[2];

        ub = (d[1] >= d[0]) ? d[1] : d[0];
    end

endmodule